library verilog;
use verilog.vl_types.all;
entity Not1bit is
    port(
        a               : in     vl_logic;
        \out\           : out    vl_logic
    );
end Not1bit;
