library verilog;
use verilog.vl_types.all;
entity Fib_TB is
end Fib_TB;
